package bus_trans_pkg;

	`include "bus_trans.SV";
	`include "derived_trans.sv";
	
endpackage : bus_trans_pkg
