

package bus_trans_v2_pkg;

	typedef enum {READ, WRITE} kind_e;
		`include "bus_trans_v2.sv"
	`include "derived_trans_v2.sv"



endpackage : bus_trans_v2_pkg
