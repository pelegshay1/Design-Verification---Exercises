module arbiter_checker (
	input clk,    // Clock
	input reset,  // Asynchronous reset active low
	input logic req_0, req_1,
	output logic gnt_0, gnt_1
);

endmodule : arbiter_checker