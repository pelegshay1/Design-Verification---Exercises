package bus_trans_pkg;
	
	`include "derived_trans.sv";
	`include "bus_trans.SV";
	
	
endpackage : bus_trans_pkg
