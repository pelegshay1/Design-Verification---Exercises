package casting_trans_pkg;
	`include "casting_trans.sv"
	`include "derived_casting_trans.sv"
endpackage : casting_trans_pkg
